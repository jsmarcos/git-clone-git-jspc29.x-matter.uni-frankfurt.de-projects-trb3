tdc_release/trb3_periph_ADA.vhd