trb3_periph_nx2.vhd