library ieee;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

package tdc_version is

  constant TDC_VERSION             : std_logic_vector(11 downto 0) := x"163";

end;
