config_default.vhd