-----------------------------------------------------------------------------
--
-- Gray Decoder
--
-----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Gray_Decoder is
  
  generic (
    WIDTH : integer := 12);             -- Register Width

  port (
    CLK_IN     : in std_logic;
    RESET_IN   : in std_logic;
    
    -- Input
    GRAY_IN    : in  std_logic_vector(WIDTH - 1 downto 0);

    -- OUTPUT
    BINARY_OUT : out std_logic_vector(WIDTH - 1 downto 0)
    );

end Gray_Decoder;


architecture Gray_Decoder of Gray_Decoder is

  signal binary_o : std_logic_vector(WIDTH - 1 downto 0);

begin  -- Gray_Decoder

  PROC_DECODER: process (CLK_IN)
  begin
    if( rising_edge(CLK_IN) ) then
      if( RESET_IN = '1' ) then
        binary_o <= (others => '0');
      else
        binary_o(WIDTH - 1) <= GRAY_IN(WIDTH - 1);
    
        for I in (WIDTH - 2) to 0 loop
          binary_o(I) <= binary_o(I + 1) xor GRAY_IN(I);
        end loop;
      end if;
    end if;
    
  end process PROC_DECODER;

  -- Output
  BINARY_OUT <= binary_o;
    
end Gray_Decoder;
