config_125.vhd