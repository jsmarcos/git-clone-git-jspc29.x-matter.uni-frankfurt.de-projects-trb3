currentRelease/cbmtof.vhd