../../cts/source/mbs_vulom_recv.vhd