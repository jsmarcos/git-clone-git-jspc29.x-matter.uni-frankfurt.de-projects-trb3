tdc_release/trb3_periph_padiwa.vhd