trb3_periph_nx1.vhd