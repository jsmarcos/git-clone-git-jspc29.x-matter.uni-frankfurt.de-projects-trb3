trb3_periph_ADA.vhd.1.6xx