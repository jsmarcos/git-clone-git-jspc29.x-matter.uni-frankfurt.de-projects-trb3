rom_encoder/ROM_encoder_3.vhd