currentRelease/trb3_periph_gpin.vhd