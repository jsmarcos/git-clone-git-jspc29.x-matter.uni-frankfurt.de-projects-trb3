../../cts/source/mainz_a2_recv.vhd