currentRelease/trb3_periph_32PinAddOn.vhd