trb3_periph_padiwa.vhd.1.6.xx