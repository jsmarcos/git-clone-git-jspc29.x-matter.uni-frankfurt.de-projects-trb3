tdc_release/cbmtof.vhd