currentRelease/trb3_periph_padiwa.vhd