tdc_release/trb3_periph_gpin.vhd