tdc_release/trb3_periph_32PinAddOn.vhd