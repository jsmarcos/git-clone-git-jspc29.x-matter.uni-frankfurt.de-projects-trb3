currentRelease/trb3_periph_ADA.vhd