trb3_components_1-6-x.vhd