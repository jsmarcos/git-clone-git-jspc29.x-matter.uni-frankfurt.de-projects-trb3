cbmtof.vhd.1.6xx