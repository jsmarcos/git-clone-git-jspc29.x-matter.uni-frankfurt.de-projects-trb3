trb3_periph_nxyter_nx1.vhd