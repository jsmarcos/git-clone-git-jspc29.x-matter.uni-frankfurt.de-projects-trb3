trb3_periph_32PinAddOn.vhd.1.6.xx